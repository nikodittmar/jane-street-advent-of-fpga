`include "control_sel.vh" 

module fpu (
    input [1:0] sel,
    input [31:0] op1,
    input [31:0] op2,
    input [31:0] op3,
    output [31:0] res
);


endmodule