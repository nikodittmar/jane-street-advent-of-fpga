module if_control (
    input br_mispred,
    input target_taken,
    input stall,
    output [1:0] pc_sel
);

endmodule