// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
`define RF_PATH   cpu.id_stage.reg_file
`define FPRF_PATH cpu.id_stage.fprf
`define DMEM_PATH cpu.mem_stage.dmem
`define IMEM_PATH cpu.imem
`define BIOS_PATH cpu.bios_mem
`define CSR_PATH  cpu.ex_stage.tohost_csr
