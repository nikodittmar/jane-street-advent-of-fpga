// List of RISC-V immediates
// Use `include "imm.vh" to use these

`ifndef IMM
`define IMM

// I-type immediates
`define IMM_I 3'b000

// S-type immediates
`define IMM_S 3'b001

// B-type immediates
`define IMM_B 3'b010

// U-type immediates
`define IMM_U 3'b011

// J-type immediates
`define IMM_J 3'b100

`endif //IMM
