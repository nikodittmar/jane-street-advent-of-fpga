`include "control_sel.vh"

module id_stage (
    input clk,
    input rst,
    input ex_flush,
    input [31:0] id_pc,
    input [31:0] id_bios_inst,
    input [31:0] id_imem_inst,
    input wb_regwen,
    input wb_fpregwen,
    input [31:0] wb_wdata,
    input [31:0] wb_inst,
    input ex_stall,
    
    output [31:0] id_target, // Branch predictor/target generator output
    output id_target_taken, // Use output of branch predictor/target generator flag
    output ex_br_taken, // Branch predictor branch taken flag
    output [31:0] ex_pc,
    output [31:0] ex_rd1,
    output [31:0] ex_rd2,
    output [31:0] ex_fd1,
    output [31:0] ex_fd2,
    output [31:0] ex_fd3,
    output [31:0] ex_imm,
    output [31:0] ex_inst,
    output id_stall
);
    wire id_reg_rst;
    wire id_reg_we;

    assign id_reg_we = ~id_stall & ~ex_stall;
    assign id_reg_rst = id_stall | ex_flush | rst;

    // MARK: InstSel

    wire [31:0] id_inst;

    wire [$clog2(`INST_SEL_NUM_INPUTS)-1:0] inst_sel = id_pc[30];
    wire [`INST_SEL_NUM_INPUTS*32-1:0] inst_mux_in;

    assign inst_mux_in[`INST_BIOS * 32 +: 32] = id_bios_inst;
    assign inst_mux_in[`INST_IMEM * 32 +: 32] = id_imem_inst;

    mux #(
        .NUM_INPUTS(`INST_SEL_NUM_INPUTS)
    ) inst_mux (
        .in(inst_mux_in),
        .sel(inst_sel),

        .out(id_inst)
    );

    // MARK: RegFile

    wire [4:0] ra1 = id_inst[19:15];
    wire [4:0] ra2 = id_inst[24:20];
    wire [4:0] wa = wb_inst[11:7];
    wire [31:0] rd1;
    wire [31:0] rd2;

    reg_file reg_file (
        .clk(clk),
        .we(wb_regwen),
        .ra1(ra1), .ra2(ra2), .wa(wa),
        .wd(wb_wdata),

        .rd1(rd1), .rd2(rd2)
    );

    // MARK: Floating Point RegFile

    wire [4:0] ra3 = id_inst[31:27];
    wire [31:0] fd1;
    wire [31:0] fd2;
    wire [31:0] fd3;

    fp_reg_file fp_reg_file (
        .clk(clk),
        .we(wb_fpregwen),
        .ra1(ra1), .ra2(ra2), .ra3(ra3), .wa(wa),
        .wd(wb_wdata),

        .rd1(fd1), .rd2(fd2), .rd3(fd3)
    );

    // MARK: ImmGen

    wire [2:0] imm_sel;
    wire [31:0] imm;

    imm_gen imm_gen (
        .inst(id_inst),
        .sel(imm_sel),

        .imm(imm)
    );

    // MARK: TargetGen
    
    wire target_gen_sel;
    wire target_gen_en;
    wire br_taken;
    
    target_gen target_gen (
        .pc(id_pc),
        .sel(target_gen_sel),
        .en(target_gen_en),
        .imm(imm),

        .target(id_target),
        .target_taken(id_target_taken),
        .branch_taken(br_taken)
    );

    // MARK: Control

    id_control control (
        .inst(id_inst),
        .ex_inst(ex_inst),
    
        .imm_sel(imm_sel),
        .target_gen_sel(target_gen_sel),
        .target_gen_en(target_gen_en),
        .stall(id_stall)
    );

    // MARK: Pipeline registers

    pipeline_reg pc_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(id_pc),

        .out(ex_pc)
    );

    pipeline_reg rd1_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(rd1),

        .out(ex_rd1)
    );

    pipeline_reg rd2_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(rd2),

        .out(ex_rd2)
    );

    pipeline_reg fd1_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(fd1),

        .out(ex_fd1)
    );

    pipeline_reg fd2_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(fd2),

        .out(ex_fd2)
    );

    pipeline_reg fd3_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(fd3),

        .out(ex_fd3)
    );

    pipeline_reg imm_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(imm),

        .out(ex_imm)
    );

    pipeline_reg #(
        .WIDTH(1)
    ) br_taken_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(br_taken),

        .out(ex_br_taken)
    );

    pipeline_reg #(
        .RESET_VAL(`NOP)
    ) inst_reg (
        .clk(clk),
        .rst(id_reg_rst),
        .we(id_reg_we),
        .in(id_inst),

        .out(ex_inst)
    );

    /*
    // System Verilog Assertions

    x_zero_is_always_zero:
        assert property ( @(posedge clk)
            (ra1 == 5'b0) |-> (rd1 == 32'b0) && (ra2 == 5'b0) |-> (rd2 == 32'b0)
        ) else $error("reading from x0 must always be zero!");
    */
    /*
    // MARK: Hazard Analysis

    reg [31:0] stall_cnt;
    
    always @(posedge clk) begin 
        if (rst) begin 
                stall_cnt <= 32'b0;
        end else begin 
            if (id_stall) begin 
                stall_cnt <= stall_cnt + 32'd1;
            end
        end
    end
    */
endmodule