`include "control_sel.vh"

module if_control (
    input rst,
    input [31:0] pc,
    input redirect_pc,
    input target_taken,
    input id_stall,
    input ex_stall,
    input flush,
    
    output reg [1:0] next_pc_sel,
    output reg [1:0] override_pc_sel,
    output reg bios_en
);

    always @(*) begin
        next_pc_sel = `PC_4;
        override_pc_sel = `PC_4;

        if (rst) begin 
            next_pc_sel = `PC_4;
            override_pc_sel = `PC_4;
        end else if (flush) begin 
            override_pc_sel = `PC_ALU;
        end else if (id_stall | ex_stall) begin 
            if (redirect_pc) begin
                next_pc_sel = `PC_ALU;
            end else if (target_taken) begin 
                next_pc_sel = `PC_TGT;
            end
        end else begin 
            if (redirect_pc) begin
                override_pc_sel = `PC_ALU;
            end else if (target_taken) begin 
                override_pc_sel = `PC_TGT;
            end
        end

        bios_en = pc[30] == `INST_BIOS;
    end

endmodule