module lzc32 (
    input  [31:0] in,
    output [5:0]  count
);
    assign count =
    (in[31]) ? 6'd0  :
    (in[30]) ? 6'd1  :
    (in[29]) ? 6'd2  :
    (in[28]) ? 6'd3  :
    (in[27]) ? 6'd4  :
    (in[26]) ? 6'd5  :
    (in[25]) ? 6'd6  :
    (in[24]) ? 6'd7  :
    (in[23]) ? 6'd8  :
    (in[22]) ? 6'd9  :
    (in[21]) ? 6'd10 :
    (in[20]) ? 6'd11 :
    (in[19]) ? 6'd12 :
    (in[18]) ? 6'd13 :
    (in[17]) ? 6'd14 :
    (in[16]) ? 6'd15 :
    (in[15]) ? 6'd16 :
    (in[14]) ? 6'd17 :
    (in[13]) ? 6'd18 :
    (in[12]) ? 6'd19 :
    (in[11]) ? 6'd20 :
    (in[10]) ? 6'd21 :
    (in[9])  ? 6'd22 :
    (in[8])  ? 6'd23 :
    (in[7])  ? 6'd24 :
    (in[6])  ? 6'd25 :
    (in[5])  ? 6'd26 :
    (in[4])  ? 6'd27 :
    (in[3])  ? 6'd28 :
    (in[2])  ? 6'd29 :
    (in[1])  ? 6'd30 :
    (in[0])  ? 6'd31 : 6'd32;
endmodule
