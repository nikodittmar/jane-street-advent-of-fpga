module if_control (
    input br_mispred,
    input target_taken,
    output [1:0] pc_sel
);

endmodule