module mem_mask (
    input [31:0] din,
    input [3:0] mask,
    output [31:0] dout
);

endmodule